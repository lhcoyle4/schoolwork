module program_counter();

endmodule