module program_terminal();
	
endmodule