module instruction_decoder();

endmodule