module uart();

endmodule