module status_register();

endmodule